library IEEE;
USE IEEE.std_logic_1164.ALL;

entity tan_lut is
port (  clk  : IN STD_LOGIC;
  deg_in: in std_logic_vector(31 downto 0);
  tan_out: out std_logic_vector(31 downto 0)
 );
end tan_lut;

ARCHITECTURE behavioral OF tan_lut IS
signal deg: std_logic_vector(7 downto 0) := deg_in(31 downto 24);
BEGIN
 tangent : PROCESS(deg)
  BEGIN
   CASE deg IS
    when "00000000" => tan_out <= "00000000000000000000000000000000"; --tan(0)
    when "00000001" => tan_out <= "00000000000001000111101011100000"; --tan(1)
    when "00000010" => tan_out <= "00000000000010001110111100110000"; --tan(2)
    when "00000011" => tan_out <= "00000000000011010110101000010000"; --tan(3)
    when "00000100" => tan_out <= "00000000000100011110010011110000"; --tan(4)
    when "00000101" => tan_out <= "00000000000101100110011001100000"; --tan(5)
    when "00000110" => tan_out <= "00000000000110101110011111010000"; --tan(6)
    when "00000111" => tan_out <= "00000000000111110110111111010000"; --tan(7)
    when "00001000" => tan_out <= "00000000001000111111011111010000"; --tan(8)
    when "00001001" => tan_out <= "00000000001010001000110011100000"; --tan(9)
    when "00001010" => tan_out <= "00000000001011010010001000000000"; --tan(10)
    when "00001011" => tan_out <= "00000000001100011100010000110000"; --tan(11)
    when "00001100" => tan_out <= "00000000001101100110110011110000"; --tan(12)
    when "00001101" => tan_out <= "00000000001110110001110001000000"; --tan(13)
    when "00001110" => tan_out <= "00000000001111111101001000100000"; --tan(14)
    when "00001111" => tan_out <= "00000000010001001001010100100000"; --tan(15)
    when "00010000" => tan_out <= "00000000010010010110010100110000"; --tan(16)
    when "00010001" => tan_out <= "00000000010011100100001001100000"; --tan(17)
    when "00010010" => tan_out <= "00000000010100110010110010100000"; --tan(18)
    when "00010011" => tan_out <= "00000000010110000010010000010000"; --tan(19)
    when "00010100" => tan_out <= "00000000010111010010111100100000"; --tan(20)
    when "00010101" => tan_out <= "00000000011000100100011101000000"; --tan(21)
    when "00010110" => tan_out <= "00000000011001110110110010010000"; --tan(22)
    when "00010111" => tan_out <= "00000000011011001010110000010000"; --tan(23)
    when "00011000" => tan_out <= "00000000011100011111100010100000"; --tan(24)
    when "00011001" => tan_out <= "00000000011101110101111101110000"; --tan(25)
    when "00011010" => tan_out <= "00000000011111001101100111110000"; --tan(26)
    when "00011011" => tan_out <= "00000000100000100110111010010000"; --tan(27)
    when "00011100" => tan_out <= "00000000100010000001110110000000"; --tan(28)
    when "00011101" => tan_out <= "00000000100011011110011010100000"; --tan(29)
    when "00011110" => tan_out <= "00000000100100111101000010000000"; --tan(30)
    when "00011111" => tan_out <= "00000000100110011101010010010000"; --tan(31)
    when "00100000" => tan_out <= "00000000100111111111100101110000"; --tan(32)
    when "00100001" => tan_out <= "00000000101001100011111100010000"; --tan(33)
    when "00100010" => tan_out <= "00000000101011001010110000010000"; --tan(34)
    when "00100011" => tan_out <= "00000000101100110100000001010000"; --tan(35)
    when "00100100" => tan_out <= "00000000101110011111101111100000"; --tan(36)
    when "00100101" => tan_out <= "00000000110000001110101111110000"; --tan(37)
    when "00100110" => tan_out <= "00000000110010000000001101000000"; --tan(38)
    when "00100111" => tan_out <= "00000000110011110100111100010000"; --tan(39)
    when "00101000" => tan_out <= "00000000110101101100111101000000"; --tan(40)
    when "00101001" => tan_out <= "00000000110111101000101001110000"; --tan(41)
    when "00101010" => tan_out <= "00000000111001101000000010100000"; --tan(42)
    when "00101011" => tan_out <= "00000000111011101011100001010000"; --tan(43)
    when "00101100" => tan_out <= "00000000111101110011100000100000"; --tan(44)
    when "00101101" => tan_out <= "00000001000000000000000000000000"; --tan(45)
    when "00101110" => tan_out <= "00000001000010010001011010000000"; --tan(46)
    when "00101111" => tan_out <= "00000001000100101000100011010000"; --tan(47)
    when "00110000" => tan_out <= "00000001000111000101000001010000"; --tan(48)
    when "00110001" => tan_out <= "00000001001001101000000010100000"; --tan(49)
    when "00110010" => tan_out <= "00000001001100010001100111010000"; --tan(50)
    when "00110011" => tan_out <= "00000001001111000010001001110000"; --tan(51)
    when "00110100" => tan_out <= "00000001010001111010011110000000"; --tan(52)
    when "00110101" => tan_out <= "00000001010100111011011001000000"; --tan(53)
    when "00110110" => tan_out <= "00000001011000000101101111000000"; --tan(54)
    when "00110111" => tan_out <= "00000001011011011001011111110000"; --tan(55)
    when "00111000" => tan_out <= "00000001011110111000101110110000"; --tan(56)
    when "00111001" => tan_out <= "00000001100010100011011011100000"; --tan(57)
    when "00111010" => tan_out <= "00000001100110011010110101000000"; --tan(58)
    when "00111011" => tan_out <= "00000001101010100000111110010000"; --tan(59)
    when "00111100" => tan_out <= "00000001101110110110101011100000"; --tan(60)
    when "00111101" => tan_out <= "00000001110011011101001011110000"; --tan(61)
    when "00111110" => tan_out <= "00000001111000010111010110010000"; --tan(62)
    when "00111111" => tan_out <= "00000001111101100110110011110000"; --tan(63)
    when "01000000" => tan_out <= "00000010000011001110000001110000"; --tan(64)
    when "01000001" => tan_out <= "00000010001001001111110111110000"; --tan(65)
    when "01000010" => tan_out <= "00000010001111101111100111100000"; --tan(66)
    when "01000011" => tan_out <= "00000010010110110001110001000000"; --tan(67)
    when "01000100" => tan_out <= "00000010011110011010000000100000"; --tan(68)
    when "01000101" => tan_out <= "00000010100110101110011111010000"; --tan(69)
    when "01000110" => tan_out <= "00000010101111110101110000110000"; --tan(70)
    when "01000111" => tan_out <= "00000010111001110111100110100000"; --tan(71)
    when "01001000" => tan_out <= "00000011000100111110010000100000"; --tan(72)
    when "01001001" => tan_out <= "00000011010001010101100110110000"; --tan(73)
    when "01001010" => tan_out <= "00000011011111001100011001000000"; --tan(74)
    when "01001011" => tan_out <= "00000011101110110110101011100000"; --tan(75)
    when "01001100" => tan_out <= "00000100000000101100001111010000"; --tan(76)
    when "01001101" => tan_out <= "00000100010101001101110100110000"; --tan(77)
    when "01001110" => tan_out <= "00000100101101000110000010110000"; --tan(78)
    when "01001111" => tan_out <= "00000101001001010000010010000000"; --tan(79)
    when "01010000" => tan_out <= "00000101101010111101101001010000"; --tan(80)
    when "01010001" => tan_out <= "00000110010100000101010100110000"; --tan(81)
    when "01010010" => tan_out <= "00000111000111011000101011100000"; --tan(82)
    when "01010011" => tan_out <= "00001000001001001111000011100000"; --tan(83)
    when "01010100" => tan_out <= "00001001100000111010111110110000"; --tan(84)
    when "01010101" => tan_out <= "00001011011011100001101100010000"; --tan(85)
    when "01010110" => tan_out <= "00001110010011001111101010110000"; --tan(86)
    when "01010111" => tan_out <= "00010011000101001100001100000000"; --tan(87)
    when "01011000" => tan_out <= "00011100101000101110010010010000"; --tan(88)
    when "01011001" => tan_out <= "00111001010010100011110101110000"; --tan(89)
    when "01011010" => tan_out <= "11111111111111111111111111111111"; --tan(90)
    when others => tan_out <= "00000000000000000000000000000000"; --tan(>90)
   end case;
  end process;
end behavioral;